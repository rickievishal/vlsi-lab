module ex1(a,b,y);
  input a,b;
  output y;
  or a1(y,a,b);
endmodule